module menu

import gg
import gx

// Menu is the menu that is drawn on the title screen.
pub struct Menu {
__global:
	x              int
	y              int
	menu_items     []MenuItem
	text_alignment TextAlignment
	selected       SelectedMenuItem
	text_color     gx.Color = gx.rgb(0xba, 0xba, 0xba)
	font_size      int      = 40
}

// Menu.new creates a new `Menu` at the given position with the given menu items.
[inline]
pub fn Menu.new(menu_items ...MenuItem) Menu {
	return Menu{
		menu_items: menu_items
	}
}

// center centers the menu relative to the window size.
pub fn (mut menu Menu) center(mut g gg.Context) {
	menu.x = g.width / 2 - menu.width(mut g) / 2
	menu.y = g.height / 2 - menu.height(mut g) / 2
}

// event handles events for the menu.
pub fn (mut menu Menu) event(event &gg.Event) {
	match event.typ {
		.key_down {
			match event.key_code {
				.up {
					menu.selected.index = (menu.selected.index - 1) % menu.menu_items.len
				}
				.down {
					menu.selected.index = (menu.selected.index + 1) % menu.menu_items.len
				}
				.left {
					mut menu_item := menu.menu_items[menu.selected.index]
					match mut menu_item {
						CycleMenuItem {
							if menu_item.selected_value > 0 {
								menu_item.cycle_left()
							}
						}
						else {}
					}
				}
				.right {
					mut menu_item := menu.menu_items[menu.selected.index]
					match mut menu_item {
						CycleMenuItem {
							if menu_item.selected_value < menu_item.values.len - 1 {
								menu_item.cycle_right()
							}
						}
						else {}
					}
				}
				.enter {
					mut menu_item := menu.menu_items[menu.selected.index]
					match mut menu_item {
						ButtonMenuItem {
							if click_fn := menu_item.on.click {
								click_fn()
							}
						}
						CycleMenuItem {
							menu_item.current_value = menu_item.selected_value
							if click_fn := menu_item.on.click {
								click_fn(menu_item.value())
							}
						}
						ToggleMenuItem {
							menu_item.toggled_on = !menu_item.toggled_on
							if toggle_fn := menu_item.on.toggle {
								toggle_fn(menu_item.toggled_on)
							} else {
								if menu_item.toggled_on {
									if toggle_on_fn := menu_item.on.toggle_on {
										toggle_on_fn()
									}
								} else {
									if toggle_off_fn := menu_item.on.toggle_off {
										toggle_off_fn()
									}
								}
							}
						}
					}
				}
				else {}
			}
		}
		else {}
	}
}

// current_item returns the currently selected menu item.
[inline]
pub fn (mut menu Menu) current_item() MenuItem {
	return menu.menu_items[menu.selected.index]
}

// width returns the width of the menu.
pub fn (mut menu Menu) width(mut g gg.Context) int {
	mut max_width := 0
	for mut menu_item in menu.menu_items {
		match mut menu_item {
			ButtonMenuItem {
				width := g.text_width(menu_item.label) + menu_item.padding.left +
					menu_item.padding.right + menu_item.border.size * 2
				if width > max_width {
					max_width = width
				}
			}
			CycleMenuItem {
				// +2 for the arrow characters and +2 for the space between
				// the arrow characters and the label.
				width := g.text_width(menu_item.label) + menu_item.padding.left +
					menu_item.padding.right + 4
				if width > max_width {
					max_width = width
				}
			}
			ToggleMenuItem {
				width := g.text_width(menu_item.text()) + menu_item.padding.left +
					menu_item.padding.right
				if width > max_width {
					max_width = width
				}
			}
		}
	}
	return max_width
}

// height returns the height of the menu.
pub fn (mut menu Menu) height(mut g gg.Context) int {
	mut height := 0
	for mut menu_item in menu.menu_items {
		match mut menu_item {
			ButtonMenuItem {
				height += g.text_height(menu_item.label) + menu_item.padding.top +
					menu_item.padding.bottom + (menu_item.border.size * 2)
			}
			CycleMenuItem {
				height += g.text_height(menu_item.label) + menu_item.padding.top +
					menu_item.padding.bottom
			}
			ToggleMenuItem {
				height += g.text_height(menu_item.text()) + menu_item.padding.top +
					menu_item.padding.bottom
			}
		}
	}
	return height
}

// draw draws the menu to the screen.
[direct_array_access]
pub fn (mut menu Menu) draw(mut g gg.Context) {
	mut offset_y := 0
	for i, mut menu_item in menu.menu_items {
		is_selected_item := i == menu.selected.index
		menu_item_color := if is_selected_item {
			menu.selected.text_color
		} else {
			menu.text_color
		}
		match mut menu_item {
			ButtonMenuItem {
				border_x := menu.x
				border_y := menu.y + offset_y
				local_offset_x := menu_item.padding.left + menu_item.border.size
				local_offset_y := menu_item.padding.top + menu_item.border.size
				button_x := menu.x + local_offset_x
				button_y := menu.y + offset_y + local_offset_y
				border_width := g.text_width(menu_item.label) + menu_item.padding.left +
					menu_item.padding.right + (menu_item.border.size * 2)
				border_height := g.text_height(menu_item.label) + menu_item.padding.top +
					menu_item.padding.bottom + (menu_item.border.size * 2)
				offset_y += border_height
				g.draw_text(button_x, button_y, menu_item.label,
					size: menu.font_size
					color: menu_item_color
				)
				if menu_item.border.size > 0 {
					g.draw_rounded_rect_empty(border_x, border_y, border_width, border_height,
						menu_item.border.radius, menu_item.border.color)
				}
				annotation_margin := 10
				if menu.selected.annotation[0].len > 0 && is_selected_item {
					annotation_width := g.text_width(menu.selected.annotation[0])
					g.draw_text(border_x - annotation_margin - annotation_width, border_y +
						local_offset_y, menu.selected.annotation[0],
						size: menu.font_size
						color: menu.selected.text_color
					)
				}
				if menu.selected.annotation[1].len > 0 && is_selected_item {
					g.draw_text(border_x + border_width + annotation_margin, border_y +
						local_offset_y, menu.selected.annotation[1],
						size: menu.font_size
						color: menu.selected.text_color
					)
				}
			}
			CycleMenuItem {
				local_offset_x := menu_item.padding.left
				local_offset_y := menu_item.padding.top
				cycle_x := menu.x + local_offset_x
				cycle_y := menu.y + offset_y + local_offset_y
				offset_y += g.text_height(menu_item.label) + menu_item.padding.top +
					menu_item.padding.bottom

				value_color := if menu_item.selected_value == menu_item.current_value {
					menu.text_color
				} else {
					gx.rgb(0xca, 0x33, 0x5a)
				}
				label := '${menu_item.label}: '
				cycle_left := '< '
				cycle_right := ' >'
				value := menu_item.value()
				is_first_item := menu_item.selected_value == 0
				is_last_item := menu_item.selected_value == menu_item.values.len - 1
				g.draw_text(cycle_x, cycle_y, label,
					size: menu.font_size
					color: menu_item_color
				)
				g.draw_text(cycle_x + g.text_width(label), cycle_y, cycle_left,
					size: menu.font_size
					color: if is_first_item {
						menu.text_color
					} else {
						menu.selected.text_color
					}
				)
				g.draw_text(cycle_x + g.text_width(label) + g.text_width(cycle_left),
					cycle_y, value,
					size: menu.font_size
					color: value_color
				)
				g.draw_text(cycle_x + g.text_width(label) + g.text_width(cycle_left) +
					g.text_width(value), cycle_y, cycle_right,
					size: menu.font_size
					color: if is_last_item {
						menu.text_color
					} else {
						menu.selected.text_color
					}
				)
			}
			ToggleMenuItem {
				border_x := menu.x
				border_y := menu.y + offset_y
				local_offset_x := menu_item.padding.left + menu_item.border.size
				local_offset_y := menu_item.padding.top + menu_item.border.size
				toggler_x := menu.x + local_offset_x
				toggler_y := menu.y + offset_y + local_offset_y
				border_width := g.text_width(menu_item.text()) + menu_item.padding.left +
					menu_item.padding.right + (menu_item.border.size * 2)
				border_height := g.text_height(menu_item.text()) + menu_item.padding.top +
					menu_item.padding.bottom + (menu_item.border.size * 2)
				offset_y += border_height
				g.draw_text(toggler_x, toggler_y, menu_item.text(),
					size: menu.font_size
					color: menu_item_color
				)
				if menu_item.border.size > 0 {
					g.draw_rounded_rect_empty(border_x, border_y, border_width, border_height,
						menu_item.border.radius, menu_item.border.color)
				}
			}
		}
	}
}

// todo: replace with anonymous struct.
// vfmt currently has a bug that prevents this.
pub struct SelectedMenuItem {
mut:
	index      int
	text_color gx.Color = gx.white
	// annotation is the character used to denote the selected item.
	/**
	 * example if annotation[0] is '>'
	 *   > selected
	 *     unselected
	 *     unselected
	 * example if annotation[1] is '<'
	 *     unselected <
	 *     selected
	 *     unselected
	**/
	annotation [2]string
}

// TextAlignment is the alignment of the text.
pub enum TextAlignment {
	left
	right
	center
	justify
}

// Padding is the extra distance given around an item (in pixels).
pub struct Padding {
__global:
	top    int
	right  int
	bottom int
	left   int
}

// Padding.new creates a new `Padding` with the same padding on all sides.
[inline]
pub fn Padding.new(padding int) Padding {
	return Padding{padding, padding, padding, padding}
}

// Padding.yx creates a new `Padding` with the given padding on the y (top
// and bottom) and x (left and right) axes.
[inline]
pub fn Padding.yx(y int, x int) Padding {
	return Padding{y, x, y, x}
}
