module main

// Pos is a position in 2D space.
interface Pos {
mut:
	x f32
	y f32
}
