module main

import core

fn main() {
	mut game := core.Game.new()
	game.run()
}
