module core

// background textures are orderd in the way they are drawn.
const const_textures = {
	'stringstar-fields': {
		'background_0': $embed_file('../assets/stringstar-fields/background_0.png')
		'background_1': $embed_file('../assets/stringstar-fields/background_1.png')
		'background_2': $embed_file('../assets/stringstar-fields/background_2.png')
		'tileset':      $embed_file('../assets/stringstar-fields/tileset.png')
		'level':        $embed_file('../assets/stringstar-fields/example_no_background.png')
	}
}
